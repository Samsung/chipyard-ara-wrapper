// Dummy file used for source flattener.
